`include "RegisterFile.v"
module test_Register_File;
	wire [31:0]PA, PB, PC, pc_out;
	reg [31:0] PW, pc_in, pc_plus_4;
	reg [3:0] RA, RB, RC;
	wire [15:0] Registers_Enable;
	wire [31:0] R15, R14, R13, R12, R11, R10, R9, R8, R7, R6, R5, R4, R3, R2, R1, R0;
	reg [3:0] RW;
	reg  load, Clk, BL_true, pc_enable;
	
 	Register_File RF(PA, PB, PC, PW, RA, RB, RC, RW, pc_out, pc_in, pc_enable,  pc_plus_4, BL_true, load, Clk);
 	
	initial #1000 $finish;
	initial begin
	    PW = 32'b00000000000000000000000000000111;
	    RA = 4'b0011;
	    RB = 4'b1000;
	    RC = 4'b0110;
	    RW = 4'b0011;
	    pc_in = 32'b00000000000000000000000000000000;
	    pc_enable = 1'b1;
	    pc_plus_4 = 32'b00000000000000000000000000000100;
	    BL_true = 1'b0;
	    load = 1'b1;
	    Clk = 1'b0;
	    repeat(20)
	    #20 Clk <= ~Clk;
	end
	
	initial fork
	
	#20 PW = 32'b00000000001100000110000000000111;
	#20 RW = 4'b0001;
	#20 RA = 4'b0001;

	#40 PW = 32'b00111000001100000110000001111000;
	#40 RW = 4'b0010;
	#40 RB = 4'b0010;
	
	#60 PW = 32'b00000000000000000000000000000001;
	#60 RW = 4'b0011;
	#60 RC = 4'b0011;
	
	#80 PW = 32'b00111000000000000000000000000000;
	#80 RW = 4'b0100;
	#80 RA = 4'b0100;
	
	#100 PW = 32'b00000000001111000000000111100000;
	#100 RW = 4'b0101;
	#100 RB = 4'b0101;

	#120 PW = 32'b00000000000000000000000000000111;
	#120 RW = 4'b0110;
	#120 RC = 4'b0110;
	
	#140 PW = 32'b00111000000000000000000001111111;
	#140 RW = 4'b0111;
	#140 RA = 4'b0111;
	
	#160 PW = 32'b11111110000000000000000000000001;
	#160 RW = 4'b1000;
	#160 RB = 4'b1000;
	
	#180 PW = 32'b00000000000001111100000000000000;
	#180 RW = 4'b1001;
	#180 RC = 4'b1001;
	
	#200 PW = 32'b10000000000000000000000000000001;
	#200 RW = 4'b1010;
	#200 RA = 4'b1010;
	
	#220 PW = 32'b00000000001100000000000000000000;
	#220 RW = 4'b1011;
	#220 RB = 4'b1011;
	
	#240 PW = 32'b00000000000000000110000001111000;
	#240 RW = 4'b1100;
	#240 RC = 4'b1100;
	
	#260 PW = 32'b00000000000000000000000011111111;
	#260 RW = 4'b1101;
	#260 RA = 4'b1101;
	
	#280 PW = 32'b00000000000000000001111100000000;
	#280 RW = 4'b1110;
	#280 RB = 4'b1110;
	
	#300 PW = 32'b00000010101010101010101010101010;
	#300 RW = 4'b1111;
	#300 RC = 4'b1111;

	#340 PW = 32'b11111111111111110000000000000000;
	#340 RW = 4'b0001;
	#340 RB = 4'b0001;
	#340 RA = 4'b1111;	

    // #380 BL_true = 1'b1;
	#380 PW = 32'b00000000001100000110000000000111;
	#380 RB = 4'b1110;
    #380 RW = 4'b1110;
    
	join 
	initial begin
	$display("Program Counter PA PB PC RA RB RC PW RW load Clk Time");
	$monitor (" %b %b %b %b %b %b %b %b %b %b %b ", pc_out, PA, PB, PC, RA, RB, RC, PW, RW, load, Clk, $time);
    end
endmodule